.SUBCKT bufbdk Z I VSS VDD
M1 net105 net140 net106 net106 NMOS W=1.028u L=0.18u nf=1
M2 net107 net141 net108 net108 NMOS W=1.028u L=0.18u nf=1
M3 net106 net142 net107 net107 NMOS W=1.028u L=0.18u nf=1
M4 net104 net143 net105 net105 NMOS W=1.028u L=0.18u nf=1
M5 net103 net144 net104 net104 NMOS W=1.028u L=0.18u nf=1
M6 net102 net145 net103 net103 NMOS W=1.028u L=0.18u nf=1
M7 net101 net146 net102 net102 NMOS W=1.028u L=0.18u nf=1
M8 net100 net147 net101 net101 NMOS W=1.028u L=0.18u nf=1
M9 net100 net148 net99 net99 NMOS W=1.028u L=0.18u nf=1
M10 net98 net149 net99 net99 NMOS W=1.028u L=0.18u nf=1
M11 net97 net150 net98 net98 NMOS W=1.028u L=0.18u nf=1
M12 net96 net151 net97 net97 NMOS W=1.028u L=0.18u nf=1
M13 net95 net152 net96 net96 NMOS W=1.028u L=0.18u nf=1
M14 net108 net153 net109 net109 NMOS W=1.022u L=0.18u nf=1
M15 net110 net154 net95 net95 NMOS W=0.472u L=0.18u nf=1
M16 net110 net155 net111 net111 NMOS W=0.472u L=0.18u nf=1
M17 net111 net156 net112 net112 NMOS W=0.472u L=0.18u nf=1
M18 net116 net121 net83 net83 PMOS W=2.689u L=0.18u nf=1
M19 net90 net122 net91 net91 PMOS W=1.089u L=0.18u nf=1
M20 net120 net123 net90 net90 PMOS W=2.689u L=0.18u nf=1
M21 net120 net124 net89 net89 PMOS W=2.689u L=0.18u nf=1
M22 net119 net125 net89 net89 PMOS W=2.689u L=0.18u nf=1
M23 net119 net126 net88 net88 PMOS W=2.689u L=0.18u nf=1
M24 net115 net127 net88 net88 PMOS W=2.689u L=0.18u nf=1
M25 net118 net128 net87 net87 PMOS W=2.689u L=0.18u nf=1
M26 net82 net129 net83 net83 PMOS W=2.689u L=0.18u nf=1
M27 net116 net130 net84 net84 PMOS W=2.689u L=0.18u nf=1
M28 net114 net131 net84 net84 PMOS W=2.689u L=0.18u nf=1
M29 net114 net132 net85 net85 PMOS W=2.689u L=0.18u nf=1
M30 net117 net133 net86 net86 PMOS W=2.689u L=0.18u nf=1
M31 net115 net134 net87 net87 PMOS W=2.689u L=0.18u nf=1
M32 net118 net135 net86 net86 PMOS W=2.689u L=0.18u nf=1
M33 net117 net136 net85 net85 PMOS W=2.689u L=0.18u nf=1
M34 net93 net137 net94 net94 PMOS W=1.511u L=0.18u nf=1
M35 net82 net138 net92 net92 PMOS W=2.228u L=0.18u nf=1
M36 net92 net139 net93 net93 PMOS W=1.389u L=0.18u nf=1
.ends bufbdk