.SUBCKT	an02d7	Z	A1	A2	VDD	VSS
M1	U3_drain	A2	VDD	VDD	P	L=0.184U	W=1.86U	
+	PD=.820U
M2	U3_drain	A1	VDD	VDD	P	L=0.184U	W=1.86U	
+	PD=.820U
M3	Z	U3_drain	VDD	VDD	P	L=0.185167U	W=14.37U	
+	PD=1.505U
M4	u2_drain	A2	VSS	VSS	N	L=0.18U	W=1.01U	
+	PD=.700U
M5	U3_drain	A1	u2_drain	VSS	N	L=0.188U	W=1.01U	
+	PS=.700U	PD=.700U
M6	Z	U3_drain	VSS	VSS	N	L=0.18U	W=5.05U	
+	PD=1.382U

.ENDS	an02d7

.SUBCKT	bufbdk	Z	I	VDD	VSS
M1	Z	U2_gate	VDD	VDD	P	L=0.182812U	W=40.68U
M2	U2_gate	I	VDD	VDD	P	L=0.183333U	W=5.03U
M3	Z	U2_gate	VSS	VSS	N	L=0.18U	W=14.41U
M4	U2_gate	I	VSS	VSS	N	L=0.18U	W=1.41U

.ENDS	bufbdk

.SUBCKT	invbda	ZN	I	VDD	VSS
M1	ZN	I	VSS	VSS	N	L=0.18U	W=6.98U
M2	ZN	I	VDD	VDD	P	L=0.182333U	W=20.13U

.ENDS	invbda

.SUBCKT	nr02d7	ZN	A4	A5	VDD	VSS
M1	U36_out	U36_in	VSS	VSS	N	L=0.18U	W=0.97U	
M2	U36_out	U36_in	VDD	VDD	P	L=0.183U	W=2.26U	
M3	ZN	U36_out	VSS	VSS	N	L=0.1865U	W=5.05U	
M4	ZN11	U36_out	VDD	VDD	P	L=0.18U	W=14.34U	
M5	U36_in	A4	VSS	VSS	N	L=0.18U	W=0.42U	
M6	U36_in	A2	VSS	VSS	N	L=0.18U	W=0.42U	
M7	U36_in	A2	u1_source	VDD	P	L=0.187U	W=2.12U	
M8	VDD	A1	u1_source	VDD	P	L=0.183U	W=2.12U	

.ENDS	nr02d7
